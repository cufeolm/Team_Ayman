`include "GUVM_sequence.sv"
`include "child_sequence.sv"
`include "python_sequence.sv"
`include"add_seq.sv"
`include"bief_seq.sv"
`include"subcc_seq.sv"
`include"load_double_seq.sv"
