`include "GUVM_sequence.sv"
`include"add_seq.sv"
