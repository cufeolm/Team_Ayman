`include "add.svh"
`include "test.svh"
`include "jal.svh"
`include "load.svh"
`include "store.svh"
`include "nop.svh"
`include "addcc.svh"
`include "addx.svh"
`include "addxcc.svh"
`include "bief.svh"
`include "bier.svh"
`include "bvsf.svh"
`include "bcsf.svh"
`include "bnegf.svh"
`include "ba.svh"
`include "jalr.svh"
`include "jalr_cpc.svh"
`include "jalrr.svh"
`include "subcc.svh"
`include "bigtoer.svh"
`include "biltr.svh"
`include "bigtoeru.svh"
`include "biltru.svh"
`include "lwrr.svh"
`include "lsbma.svh"
`include "lshma.svh"
`include "lubma.svh"
`include "luhma.svh"
`include "lwma.svh"
`include "lw.svh"
`include "lsbmarr.svh" // riscy extension instruction
`include "lshmarr.svh" // riscy extension instruction
`include "lubmarr.svh" // riscy extension instruction
`include "luhmarr.svh" // riscy extension instruction
`include "lwmarr.svh" // riscy extension instruction
`include "ldd.svh"
`include "lddrr.svh"
`include"rdpsr.svh"
`include "sbma.svh"
`include "shma.svh"
`include "swma.svh"
