`include "add.svh"
`include "test.svh"
`include "jal.svh"
`include "load.svh"
`include "store.svh"
`include "nop.svh"
`include "addcc.svh"
`include "addx.svh"
`include "bief.svh"
`include "bvsf.svh"
`include "bcsf.svh"
`include "bnegf.svh"
`include "ba.svh"
`include "jalr.svh"
`include "jalr_cpc.svh"
`include "jalrr.svh"
`include "subcc.svh"