`include "GUVM_test.sv"
`include"add_test.sv"